module  display7seg(dp, dado, leds);
input dp;
input [3:0] dado;
output reg [7:0] leds;
endmodule